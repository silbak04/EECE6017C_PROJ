`define     BCD_0       4'h0
`define     BCD_1       4'h1
`define     BCD_2       4'h2
`define     BCD_3       4'h3
`define     BCD_4       4'h4
`define     BCD_5       4'h5
`define     BCD_6       4'h6
`define     BCD_7       4'h7
`define     BCD_8       4'h8
`define     BCD_9       4'h9
`define     BCD_A       4'hA
`define     BCD_B       4'hB
`define     BCD_C       4'hC
`define     BCD_D       4'hD
`define     BCD_E       4'hE
`define     BCD_BLANK   4'hF

// vim: set filetype=verilog: 
