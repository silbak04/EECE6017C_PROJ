`include "constants.vh"

/*--==========================================================================--*/
//--================================= VERILOG ==================================--
//--============================================================================--
//--                                                                            --
//-- FILE NAME: top.v                                                           --
//--                                                                            --
//-- DATE: 9/30/2012                                                            --
//--                                                                            --
//-- DESIGNER: Samir Silbak                                                     --
//--                                                                            --
//-- DESCRIPTION: top                                                           --
//--                                                                            --
//--============================================================================--
//--================================= VERILOG ==================================--
/*--===========================================================================--*/

module top (
    input CLOCK_50,

    input [3:0] KEY,
    input [9:0] SW,

    output [7:0] LEDG,
    output [9:0] LEDR,

    output [6:0] HEX0,
    output [6:0] HEX1,
    output [6:0] HEX2,
    output [6:0] HEX3
);

/*--============================================================--*/
/*--                        KEY MAPPINGS                        --*/
/*--============================================================--*/

    assign clk = CLOCK_50;
    assign rst = ~(KEY[0]);

    assign start = ~(KEY[3]);
    
/*--============================================================--*/
/*--                      START/STOP PROGRAM                    --*/
/*--============================================================--*/

    reg run = 0;
    reg stop = 0;

    always @ (posedge start, posedge rst) begin
        if (rst) begin
            run = 0;
            stop = 0;
        end else begin
            run = ~run;
            if (run == 0) stop = 1;
            else stop = 0;
        end
    end

    assign LEDG[7] = run;
    assign LEDG[6] = stop;

/*--============================================================--*/
/*--                    RANDOM NUMBER GENERATOR                 --*/
/*--============================================================--*/

    wire [7:0] rand_num;

    rng rng (
        .clk(clk),
        .en(run),
        .rst(rst),
        .out(rand_num)
    );

/*--============================================================--*/
/*--                        DIVIDE BY THREE                     --*/
/*--============================================================--*/

    wire [7:0] div_num;

    divide_by_three divider1 (
        .dividend(rand_num),
        .quotient(div_num)
    );

/*--============================================================--*/
/*--                          SUM THREE                         --*/
/*--============================================================--*/

    wire [7:0] sum_val;

    sum_3 sum_3 (
        .clk(clk),
        .rst(rst),
        .en(run),
        .in(div_num),
        .out(sum_val)
    );

    assign LEDR [7:0] = sum_val;

/*--============================================================--*/
/*--                          COUNTER                           --*/
/*--============================================================--*/

    counter counter (
        .clk(clk),
        .rst(rst),
        .en(run),
        .stop(stop),

        .sev_seg0(HEX0),
        .sev_seg1(HEX1),
        .sev_seg2(HEX2),
        .sev_seg3(HEX3)
    );

endmodule
