`define OFF                 4'hA
`define NEGATIVE            4'hB

// vim: set filetype=verilog: 
