`define     BCD_0       4'h00
`define     BCD_1       4'h01
`define     BCD_2       4'h02
`define     BCD_3       4'h03
`define     BCD_4       4'h04
`define     BCD_5       4'h05
`define     BCD_6       4'h06
`define     BCD_7       4'h07
`define     BCD_8       4'h08
`define     BCD_9       4'h09
`define     BCD_A       4'h0A
`define     BCD_B       4'h0B
`define     BCD_C       4'h0C
`define     BCD_D       4'h0D
`define     BCD_E       4'h0E
`define     BCD_BLANK   4'h0F

// vim: set filetype=verilog: 
