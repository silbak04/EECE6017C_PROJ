`define OFF                 4'hA
`define NEGATIVE            4'hB
/*`define NORMAL              
`define BORDER
`define WARNING
`define EMERGENCY*/

// vim: set filetype=verilog: 
