/*--==========================================================================--*/
//--================================= VERILOG ==================================--
//--============================================================================--
//--                                                                            --
//-- FILE NAME: seven_seg.v                                                     --
//--                                                                            --
//-- DATE: 9/18/2012                                                            --
//--                                                                            --
//-- DESIGNER: Samir Silbak                                                     --
//--           silbak04@gmail.com                                               --
//--                                                                            --
//-- DESCRIPTION: bcd 7-seg decoder                                             --
//--                                                                            --
//--============================================================================--
//--================================= VERILOG ==================================--
/*--===========================================================================--*/

module seven_seg (
    input [3:0] bcd,
    output reg [6:0] seg
);

    initial seg = 0;

    always @ (bcd) begin

        case (bcd)
            
            4'h0: seg <= 7'b1000000;  /* -- 0 -- */       /*   _____   */
            4'h1: seg <= 7'b1111001;  /* -- 1 -- */       /*  |  0  |  */
            4'h2: seg <= 7'b0100100;  /* -- 2 -- */       /* 5|     |1 */
            4'h3: seg <= 7'b0110000;  /* -- 3 -- */       /*  |_____|  */
            4'h4: seg <= 7'b0011001;  /* -- 4 -- */       /*  |  6  |  */
            4'h5: seg <= 7'b0010010;  /* -- 5 -- */       /* 4|     |2 */
            4'h6: seg <= 7'b0000010;  /* -- 6 -- */       /*  |_____|  */
            4'h7: seg <= 7'b1011000;  /* -- 7 -- */       /*     3     */
            4'h8: seg <= 7'b0000000;  /* -- 8 -- */
            4'h9: seg <= 7'b0010000;  /* -- 9 -- */
            4'hA: seg <= 7'b1111111;  /* -- off -- */
            4'hB: seg <= 7'b0111111;  /* -- "-" -- */
            4'hC: seg <= 7'b0001001;  /* -- H -- */
            4'hE: seg <= 7'b0000110;  /* -- E -- */
            4'hD: seg <= 7'b1000111;  /* -- L -- */
            4'hF: seg <= 7'b0001100;  /* -- P -- */

            default: seg <= 7'b1110011; /* "_|" for error */

        endcase

    end

endmodule

