`define OFF                 4'hA
`define NEGATIVE            4'hB
`define BLANK_STATE         4'h0
`define BLANK_ALARM         10'h0

// vim: set filetype=verilog: 
