`include "top_header.vh"

/*--==========================================================================--*/
//--================================= VERILOG ==================================--
//--============================================================================--
//--                                                                            --
//-- FILE NAME: clk_div.v                                                       --
//--                                                                            --
//-- DATE: 9/18/2012                                                            --
//--                                                                            --
//-- DESIGNER: Samir Silbak                                                     --
//--           silbak04@gmail.com                                               --
//--                                                                            --
//-- DESCRIPTION: divides the clock down to ~1.5Hz                              --
//--                                                                            --
//--============================================================================--
//--================================= VERILOG ==================================--
/*--===========================================================================--*/

module clk_div (
    input clk, clr,
    output clk_1
);

    /* (1/50e6) * 2**25 ~ 0.67s or ~1.5Hz */
    reg [24:0] q_out;

    always @ (posedge clk or negedge clr) begin
        if (clr)
            q_out <= 0;
        else
            q_out <= q_out + 1;
    end

    assign clk_1 = q_out[24]; 

endmodule
