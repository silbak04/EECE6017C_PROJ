include "constants.vh"

/*--==========================================================================--*/
//--================================= VERILOG ==================================--
//--============================================================================--
//--                                                                            --
//-- FILE NAME: seven_seg.v                                                     --
//--                                                                            --
//-- DATE: 9/18/2012                                                            --
//--                                                                            --
//-- DESIGNER: John Brady                                                       --
//--                                                                            --
//-- DESCRIPTION: bcd 7-seg decoder                                             --
//--                                                                            --
//--============================================================================--
//--================================= VERILOG ==================================--
/*--===========================================================================--*/

module seven_seg (
    input [3:0] bcd,
    output reg [6:0] seg
);

    initial seg = 0;

    always @ (bcd) begin
        case (bcd)
            
            `BCD_0: seg <= 7'b1000000;  /* -- 0 -- */       /*   _____   */
            `BCD_1: seg <= 7'b1111001;  /* -- 1 -- */       /*  |  0  |  */
            `BCD_2: seg <= 7'b0100100;  /* -- 2 -- */       /* 5|     |1 */
            `BCD_3: seg <= 7'b0110000;  /* -- 3 -- */       /*  |_____|  */
            `BCD_4: seg <= 7'b0011001;  /* -- 4 -- */       /*  |  6  |  */
            `BCD_5: seg <= 7'b0010010;  /* -- 5 -- */       /* 4|     |2 */
            `BCD_6: seg <= 7'b0000010;  /* -- 6 -- */       /*  |_____|  */
            `BCD_7: seg <= 7'b1011000;  /* -- 7 -- */       /*     3     */
            `BCD_8: seg <= 7'b0000000;  /* -- 8 -- */
            `BCD_9: seg <= 7'b0010000;  /* -- 9 -- */
            `BCD_A: seg <= 7'b1001000;  /* -- A -- */
            `BCD_B: seg <= 7'b0000111;  /* -- B -- */
            `BCD_C: seg <= 7'b1000110;  /* -- C -- */
            `BCD_D: seg <= 7'b0100001;  /* -- D -- */
            `BCD_E: seg <= 7'b0000110;  /* -- E -- */
            `BCD_BLANK: seg <= 7'b1111111;  /* -- BLANK -- */
            
            default: seg <= 7'b0111111; /* "-" for error */

        endcase

    end

endmodule
